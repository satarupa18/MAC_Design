module multiplier(input[3:0]a,b,output[11:0]product);
assign product = a*b;
endmodule